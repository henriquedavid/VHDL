ENTITY codificadordeteclado IS
	PORT ( a : IN BIT_VECTOR(9 DOWNTO 0);
			 o1      		 : OUT BIT_VECTOR( 3 DOWNTO 0 ));
END codificadordeteclado;

ARCHITECTURE codificador OF codificadordeteclado IS
BEGIN
	WITH a SELECT
		o1 <= 
			"0000" WHEN "1000000000",
			"0001" WHEN "0100000000",
			"0010" WHEN "0010000000",
			"0011" WHEN "0001000000",
			"0100" WHEN "0000100000",
			"0101" WHEN "0000010000",
			"0110" WHEN "0000001000",
			"0111" WHEN "0000000100",
			"1000" WHEN "0000000010",
			"1001" WHEN OTHERS;
END codificador;