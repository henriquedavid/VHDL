ENTITY trabalho3 IS

END trabalho3;

ARCHITECTURE arch OF trabalho3 IS
BEGIN

END arch;